module demux_1toN #(
    parameters N = 16
) (
    ports
);
    
endmodule